module mux4 	#(parameter WIDTH=8) 
		(input logic [WIDTH-1:0] d0, d1, d2, d3,
		input logic [1:0] s,
		output logic [WIDTH-1:0] y);
	
	always_comb
	case (s)
		0: assign y = d0;
		1: assign y = d1;
		2: assign y = d2;
		3: assign y = d3;
	endcase
endmodule
